-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Sun Mar 02 11:06:29 2014"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY oscilloscope IS 
	PORT
	(
		HSYNC :  OUT  STD_LOGIC;
		SC :  OUT  STD_LOGIC;
		VSYNC :  OUT  STD_LOGIC;
		DCLK :  OUT  STD_LOGIC;
		RAS :  OUT  STD_LOGIC;
		CAS :  OUT  STD_LOGIC;
		TRG :  OUT  STD_LOGIC;
		WE :  OUT  STD_LOGIC;
		ADDR :  OUT  STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END oscilloscope;

ARCHITECTURE bdf_type OF oscilloscope IS 

COMPONENT lpm_mux0
	PORT(data0x : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 data1x : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 data2x : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 data3x : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 sel : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 result : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_counter2
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_compare0
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare3
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare4
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare5
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 alb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare1
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare2
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 alb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_counter1
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_constant0
	PORT(		 result : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT scopevram
	PORT(clk : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 cs : IN STD_LOGIC;
		 rw : IN STD_LOGIC;
		 srt : IN STD_LOGIC;
		 RAS : OUT STD_LOGIC;
		 CAS : OUT STD_LOGIC;
		 TRG : OUT STD_LOGIC;
		 WE : OUT STD_LOGIC;
		 ACK : OUT STD_LOGIC;
		 BUSY : OUT STD_LOGIC;
		 AS : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_counter3
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_counter0
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ADDRESS :  STD_LOGIC_VECTOR(17 DOWNTO 0);
SIGNAL	RESET :  STD_LOGIC;
SIGNAL	SYS_CLK :  STD_LOGIC;
SIGNAL	SYS_COUNT :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	VRAM_CLK :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	DFF_inst39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	DFF_inst13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	DFF_inst42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;
SIGNAL	SRFF_inst3 :  STD_LOGIC;


BEGIN 
HSYNC <= DFF_inst18;
SYNTHESIZED_WIRE_4 <= '1';
SYNTHESIZED_WIRE_6 <= '1';
SYNTHESIZED_WIRE_7 <= '1';
SYNTHESIZED_WIRE_9 <= '1';
SYNTHESIZED_WIRE_13 <= '1';
SYNTHESIZED_WIRE_14 <= '1';
SYNTHESIZED_WIRE_15 <= '1';
SYNTHESIZED_WIRE_16 <= '1';
SYNTHESIZED_WIRE_18 <= '1';
SYNTHESIZED_WIRE_20 <= '1';
SYNTHESIZED_WIRE_21 <= '1';
SYNTHESIZED_WIRE_23 <= '1';
SYNTHESIZED_WIRE_24 <= '1';
SYNTHESIZED_WIRE_25 <= '1';
SYNTHESIZED_WIRE_26 <= '1';
SYNTHESIZED_WIRE_27 <= '1';
SYNTHESIZED_WIRE_35 <= '1';
SYNTHESIZED_WIRE_36 <= '1';
SYNTHESIZED_WIRE_37 <= '1';
SYNTHESIZED_WIRE_39 <= '1';



b2v_ADDR_MUX : lpm_mux0
PORT MAP(data0x => ADDRESS(8 DOWNTO 0),
		 data1x => ADDRESS(17 DOWNTO 9),
		 data2x => SYNTHESIZED_WIRE_0,
		 data3x => SYNTHESIZED_WIRE_1,
		 sel => SYNTHESIZED_WIRE_2,
		 result => ADDR);


b2v_HORIZONTAL_CNT : lpm_counter2
PORT MAP(sclr => RESET,
		 clock => VRAM_CLK,
		 q => SYNTHESIZED_WIRE_42);


b2v_inst : lpm_compare0
PORT MAP(dataa => SYNTHESIZED_WIRE_42,
		 ageb => SYNTHESIZED_WIRE_5);


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_4,SYNTHESIZED_WIRE_6)
BEGIN
IF (SYNTHESIZED_WIRE_4 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '0';
ELSIF (SYNTHESIZED_WIRE_6 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	SYNTHESIZED_WIRE_44 <= SYNTHESIZED_WIRE_5;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_7,SYNTHESIZED_WIRE_9)
BEGIN
IF (SYNTHESIZED_WIRE_7 = '0') THEN
	DFF_inst13 <= '0';
ELSIF (SYNTHESIZED_WIRE_9 = '0') THEN
	DFF_inst13 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DFF_inst13 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;


b2v_inst14 : lpm_compare3
PORT MAP(dataa => SYNTHESIZED_WIRE_43,
		 ageb => SYNTHESIZED_WIRE_19);


b2v_inst15 : lpm_compare4
PORT MAP(dataa => SYNTHESIZED_WIRE_43,
		 ageb => SYNTHESIZED_WIRE_30);


b2v_inst16 : lpm_compare5
PORT MAP(dataa => SYNTHESIZED_WIRE_43,
		 alb => SYNTHESIZED_WIRE_31);


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_13,SYNTHESIZED_WIRE_14)
BEGIN
IF (SYNTHESIZED_WIRE_13 = '0') THEN
	VRAM_CLK <= '0';
ELSIF (SYNTHESIZED_WIRE_14 = '0') THEN
	VRAM_CLK <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	VRAM_CLK <= SYS_COUNT(1);
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_15,SYNTHESIZED_WIRE_16)
BEGIN
IF (SYNTHESIZED_WIRE_15 = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_16 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DFF_inst18 <= SYNTHESIZED_WIRE_44;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_34 <= NOT(SYNTHESIZED_WIRE_45);



PROCESS(SYS_CLK,SYNTHESIZED_WIRE_18,SYNTHESIZED_WIRE_20)
BEGIN
IF (SYNTHESIZED_WIRE_18 = '0') THEN
	VSYNC <= '0';
ELSIF (SYNTHESIZED_WIRE_20 = '0') THEN
	VSYNC <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	VSYNC <= SYNTHESIZED_WIRE_19;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_21,SYNTHESIZED_WIRE_23)
BEGIN
IF (SYNTHESIZED_WIRE_21 = '0') THEN
	SC <= '0';
ELSIF (SYNTHESIZED_WIRE_23 = '0') THEN
	SC <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	SC <= SYNTHESIZED_WIRE_22;
END IF;
END PROCESS;









PROCESS(SYS_CLK,SYNTHESIZED_WIRE_24,SYNTHESIZED_WIRE_25)
BEGIN
IF (SYNTHESIZED_WIRE_24 = '0') THEN
	DCLK <= '0';
ELSIF (SYNTHESIZED_WIRE_25 = '0') THEN
	DCLK <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DCLK <= DFF_inst39;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_27,SYNTHESIZED_WIRE_26)
VARIABLE synthesized_var_for_SRFF_inst3 : STD_LOGIC;
BEGIN
IF (SYNTHESIZED_WIRE_27 = '0') THEN
	synthesized_var_for_SRFF_inst3 := '0';
ELSIF (SYNTHESIZED_WIRE_26 = '0') THEN
	synthesized_var_for_SRFF_inst3 := '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	synthesized_var_for_SRFF_inst3 := (NOT(synthesized_var_for_SRFF_inst3) AND SYNTHESIZED_WIRE_28) OR (synthesized_var_for_SRFF_inst3 AND (NOT(SYNTHESIZED_WIRE_29)));
END IF;
	SRFF_inst3 <= synthesized_var_for_SRFF_inst3;
END PROCESS;




SYNTHESIZED_WIRE_22 <= VRAM_CLK AND DFF_inst13 AND SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_32 AND SYNTHESIZED_WIRE_45;



SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_34 AND DFF_inst42;




PROCESS(SYS_CLK,SYNTHESIZED_WIRE_35,SYNTHESIZED_WIRE_36)
BEGIN
IF (SYNTHESIZED_WIRE_35 = '0') THEN
	DFF_inst39 <= '0';
ELSIF (SYNTHESIZED_WIRE_36 = '0') THEN
	DFF_inst39 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DFF_inst39 <= VRAM_CLK;
END IF;
END PROCESS;





PROCESS(SYS_CLK,SYNTHESIZED_WIRE_37,SYNTHESIZED_WIRE_39)
BEGIN
IF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst42 <= '0';
ELSIF (SYNTHESIZED_WIRE_39 = '0') THEN
	DFF_inst42 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DFF_inst42 <= SYNTHESIZED_WIRE_45;
END IF;
END PROCESS;




b2v_inst6 : lpm_compare1
PORT MAP(dataa => SYNTHESIZED_WIRE_42,
		 ageb => SYNTHESIZED_WIRE_32);


b2v_inst7 : lpm_compare2
PORT MAP(dataa => SYNTHESIZED_WIRE_42,
		 alb => SYNTHESIZED_WIRE_45);




b2v_ROW_TRANSFER_COUNTER : lpm_counter1
PORT MAP(sclr => RESET,
		 clock => DFF_inst18,
		 q => SYNTHESIZED_WIRE_0);


b2v_SRT_COL_START : lpm_constant0
PORT MAP(		 result => SYNTHESIZED_WIRE_1);


b2v_STATE_MACHINE : scopevram
PORT MAP(clk => SYS_CLK,
		 reset => RESET,
		 srt => SRFF_inst3,
		 RAS => RAS,
		 CAS => CAS,
		 TRG => TRG,
		 WE => WE,
		 ACK => SYNTHESIZED_WIRE_29,
		 AS => SYNTHESIZED_WIRE_2);


b2v_VERTICAL_CNT : lpm_counter3
PORT MAP(sclr => RESET,
		 clock => SYNTHESIZED_WIRE_44,
		 q => SYNTHESIZED_WIRE_43);


b2v_VRAM_CLOCK : lpm_counter0
PORT MAP(sclr => RESET,
		 clock => SYS_CLK,
		 q => SYS_COUNT);


END bdf_type;