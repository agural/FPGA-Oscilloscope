-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Tue Mar 04 12:57:31 2014"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY oscilloscope IS 
	PORT
	(
		RESET_IN :  IN  STD_LOGIC;
		CLK_IN :  IN  STD_LOGIC;
		HSYNC :  OUT  STD_LOGIC;
		SC :  OUT  STD_LOGIC;
		VSYNC :  OUT  STD_LOGIC;
		DCLK :  OUT  STD_LOGIC;
		SRT :  OUT  STD_LOGIC
	);
END oscilloscope;

ARCHITECTURE bdf_type OF oscilloscope IS 

COMPONENT lpm_counter2
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 cnt_en : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_compare0
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare3
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare4
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare5
	PORT(dataa : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
		 alb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare1
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 ageb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_compare2
	PORT(dataa : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 alb : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT lpm_counter3
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);
END COMPONENT;

COMPONENT lpm_counter0
	PORT(sclr : IN STD_LOGIC;
		 clock : IN STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	RESET :  STD_LOGIC;
SIGNAL	SYS_CLK :  STD_LOGIC;
SIGNAL	SYS_COUNT :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	VRAM_CLK :  STD_LOGIC;
SIGNAL	DFF_inst28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	DFF_inst42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	DFF_inst13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_3 <= '1';
SYNTHESIZED_WIRE_4 <= '1';
SYNTHESIZED_WIRE_6 <= '1';
SYNTHESIZED_WIRE_10 <= '1';
SYNTHESIZED_WIRE_11 <= '1';
SYNTHESIZED_WIRE_12 <= '1';
SYNTHESIZED_WIRE_13 <= '1';
SYNTHESIZED_WIRE_15 <= '1';
SYNTHESIZED_WIRE_17 <= '1';
SYNTHESIZED_WIRE_18 <= '1';
SYNTHESIZED_WIRE_20 <= '1';
SYNTHESIZED_WIRE_21 <= '1';
SYNTHESIZED_WIRE_22 <= '1';
SYNTHESIZED_WIRE_23 <= '1';
SYNTHESIZED_WIRE_24 <= '1';
SYNTHESIZED_WIRE_29 <= '1';
SYNTHESIZED_WIRE_30 <= '1';
SYNTHESIZED_WIRE_31 <= '1';
SYNTHESIZED_WIRE_33 <= '1';



b2v_HORIZONTAL_CNT : lpm_counter2
PORT MAP(sclr => RESET,
		 clock => VRAM_CLK,
		 cnt_en => DFF_inst28,
		 q => SYNTHESIZED_WIRE_39);


b2v_inst : lpm_compare0
PORT MAP(dataa => SYNTHESIZED_WIRE_39,
		 ageb => SYNTHESIZED_WIRE_2);


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_1,SYNTHESIZED_WIRE_3)
BEGIN
IF (SYNTHESIZED_WIRE_1 = '0') THEN
	SYNTHESIZED_WIRE_41 <= '0';
ELSIF (SYNTHESIZED_WIRE_3 = '0') THEN
	SYNTHESIZED_WIRE_41 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_2;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_4,SYNTHESIZED_WIRE_6)
BEGIN
IF (SYNTHESIZED_WIRE_4 = '0') THEN
	DFF_inst13 <= '0';
ELSIF (SYNTHESIZED_WIRE_6 = '0') THEN
	DFF_inst13 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DFF_inst13 <= SYNTHESIZED_WIRE_5;
END IF;
END PROCESS;


b2v_inst14 : lpm_compare3
PORT MAP(dataa => SYNTHESIZED_WIRE_40,
		 ageb => SYNTHESIZED_WIRE_16);


b2v_inst15 : lpm_compare4
PORT MAP(dataa => SYNTHESIZED_WIRE_40,
		 ageb => SYNTHESIZED_WIRE_34);


b2v_inst16 : lpm_compare5
PORT MAP(dataa => SYNTHESIZED_WIRE_40,
		 alb => SYNTHESIZED_WIRE_35);


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_10,SYNTHESIZED_WIRE_11)
BEGIN
IF (SYNTHESIZED_WIRE_10 = '0') THEN
	VRAM_CLK <= '0';
ELSIF (SYNTHESIZED_WIRE_11 = '0') THEN
	VRAM_CLK <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	VRAM_CLK <= SYS_COUNT(1);
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_12,SYNTHESIZED_WIRE_13)
BEGIN
IF (SYNTHESIZED_WIRE_12 = '0') THEN
	HSYNC <= '0';
ELSIF (SYNTHESIZED_WIRE_13 = '0') THEN
	HSYNC <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	HSYNC <= SYNTHESIZED_WIRE_41;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_28 <= NOT(SYNTHESIZED_WIRE_42);



PROCESS(SYS_CLK,SYNTHESIZED_WIRE_15,SYNTHESIZED_WIRE_17)
BEGIN
IF (SYNTHESIZED_WIRE_15 = '0') THEN
	VSYNC <= '0';
ELSIF (SYNTHESIZED_WIRE_17 = '0') THEN
	VSYNC <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	VSYNC <= SYNTHESIZED_WIRE_16;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_18,SYNTHESIZED_WIRE_20)
BEGIN
IF (SYNTHESIZED_WIRE_18 = '0') THEN
	SC <= '0';
ELSIF (SYNTHESIZED_WIRE_20 = '0') THEN
	SC <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	SC <= SYNTHESIZED_WIRE_19;
END IF;
END PROCESS;








PROCESS(VRAM_CLK,SYNTHESIZED_WIRE_21,SYNTHESIZED_WIRE_22)
BEGIN
IF (SYNTHESIZED_WIRE_21 = '0') THEN
	DFF_inst28 <= '0';
ELSIF (SYNTHESIZED_WIRE_22 = '0') THEN
	DFF_inst28 <= '1';
ELSIF (RISING_EDGE(VRAM_CLK)) THEN
	DFF_inst28 <= VRAM_CLK;
END IF;
END PROCESS;


PROCESS(SYS_CLK,SYNTHESIZED_WIRE_23,SYNTHESIZED_WIRE_24)
BEGIN
IF (SYNTHESIZED_WIRE_23 = '0') THEN
	DCLK <= '0';
ELSIF (SYNTHESIZED_WIRE_24 = '0') THEN
	DCLK <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	DCLK <= SYNTHESIZED_WIRE_43;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_38 <= NOT(SYNTHESIZED_WIRE_41);






SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_25 AND SYNTHESIZED_WIRE_26;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_42;


SRT <= SYNTHESIZED_WIRE_28 AND DFF_inst42;





PROCESS(SYS_CLK,SYNTHESIZED_WIRE_29,SYNTHESIZED_WIRE_30)
BEGIN
IF (SYNTHESIZED_WIRE_29 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_30 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(SYS_CLK)) THEN
	SYNTHESIZED_WIRE_43 <= VRAM_CLK;
END IF;
END PROCESS;





PROCESS(VRAM_CLK,SYNTHESIZED_WIRE_31,SYNTHESIZED_WIRE_33)
BEGIN
IF (SYNTHESIZED_WIRE_31 = '0') THEN
	DFF_inst42 <= '0';
ELSIF (SYNTHESIZED_WIRE_33 = '0') THEN
	DFF_inst42 <= '1';
ELSIF (RISING_EDGE(VRAM_CLK)) THEN
	DFF_inst42 <= SYNTHESIZED_WIRE_42;
END IF;
END PROCESS;




SYNTHESIZED_WIRE_42 <= DFF_inst13 AND SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35;


b2v_inst6 : lpm_compare1
PORT MAP(dataa => SYNTHESIZED_WIRE_39,
		 ageb => SYNTHESIZED_WIRE_25);


b2v_inst7 : lpm_compare2
PORT MAP(dataa => SYNTHESIZED_WIRE_39,
		 alb => SYNTHESIZED_WIRE_26);




b2v_VERTICAL_CNT : lpm_counter3
PORT MAP(sclr => RESET,
		 clock => SYNTHESIZED_WIRE_38,
		 q => SYNTHESIZED_WIRE_40);


b2v_VRAM_CLOCK : lpm_counter0
PORT MAP(sclr => RESET,
		 clock => SYS_CLK,
		 q => SYS_COUNT);

SYS_CLK <= CLK_IN;
RESET <= RESET_IN;

END bdf_type;