-- proc.vhd

-- Generated using ACDS version 13.1 162 at 2014.06.12.19:57:24

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity proc is
	port (
		clk_clk                                   : in    std_logic                     := '0';             --         clk.clk
		bridge_out_VRAM_ctrl_tcm_data_out         : inout std_logic_vector(15 downto 0) := (others => '0'); --  bridge_out.VRAM_ctrl_tcm_data_out
		bridge_out_VRAM_ctrl_tcm_chipselect_n_out : out   std_logic_vector(0 downto 0);                     --            .VRAM_ctrl_tcm_chipselect_n_out
		bridge_out_VRAM_ctrl_tcm_waitrequest_in   : in    std_logic_vector(0 downto 0)  := (others => '0'); --            .VRAM_ctrl_tcm_waitrequest_in
		bridge_out_data                           : inout std_logic_vector(7 downto 0)  := (others => '0'); --            .data
		bridge_out_VRAM_ctrl_tcm_address_out      : out   std_logic_vector(18 downto 0);                    --            .VRAM_ctrl_tcm_address_out
		bridge_out_r_w                            : out   std_logic_vector(0 downto 0);                     --            .r_w
		bridge_out_RAM_ctrl_tcm_chipselect_n_out  : out   std_logic_vector(0 downto 0);                     --            .RAM_ctrl_tcm_chipselect_n_out
		bridge_out_VRAM_ctrl_tcm_write_n_out      : out   std_logic_vector(0 downto 0);                     --            .VRAM_ctrl_tcm_write_n_out
		bridge_out_ROM_ctrl_tcm_chipselect_n_out  : out   std_logic_vector(0 downto 0);                     --            .ROM_ctrl_tcm_chipselect_n_out
		bridge_out_address                        : out   std_logic_vector(15 downto 0);                    --            .address
		key_input_export                          : in    std_logic_vector(19 downto 0) := (others => '0'); --   key_input.export
		adc_raw_export                            : in    std_logic_vector(23 downto 0) := (others => '0'); --     adc_raw.export
		trig_int_export                           : in    std_logic_vector(7 downto 0)  := (others => '0'); --    trig_int.export
		adc_ctrl_export                           : out   std_logic_vector(7 downto 0);                     --    adc_ctrl.export
		adc_rate_export                           : out   std_logic_vector(31 downto 0);                    --    adc_rate.export
		trig_ctrl_export                          : out   std_logic_vector(7 downto 0);                     --   trig_ctrl.export
		trig_level_export                         : out   std_logic_vector(7 downto 0);                     --  trig_level.export
		trig_delay_export                         : out   std_logic_vector(15 downto 0);                    --  trig_delay.export
		trig_errorr_export                        : out   std_logic_vector(7 downto 0);                     -- trig_errorr.export
		test_inp_export                           : in    std_logic_vector(31 downto 0) := (others => '0')  --    test_inp.export
	);
end entity proc;

architecture rtl of proc is
	component proc_PROC is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(20 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component proc_PROC;

	component proc_RAM_ctrl is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(15 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component proc_RAM_ctrl;

	component proc_ROM_ctrl is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(15 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component proc_ROM_ctrl;

	component proc_PIN_share is
		port (
			clk_clk                        : in  std_logic                     := 'X';             -- clk
			reset_reset                    : in  std_logic                     := 'X';             -- reset
			request                        : out std_logic;                                        -- request
			grant                          : in  std_logic                     := 'X';             -- grant
			VRAM_ctrl_tcm_address_out      : out std_logic_vector(18 downto 0);                    -- VRAM_ctrl_tcm_address_out_out
			VRAM_ctrl_tcm_waitrequest_in   : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- VRAM_ctrl_tcm_waitrequest_in_in
			VRAM_ctrl_tcm_write_n_out      : out std_logic_vector(0 downto 0);                     -- VRAM_ctrl_tcm_write_n_out_out
			VRAM_ctrl_tcm_data_out         : out std_logic_vector(15 downto 0);                    -- VRAM_ctrl_tcm_data_out_out
			VRAM_ctrl_tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- VRAM_ctrl_tcm_data_out_in
			VRAM_ctrl_tcm_data_outen       : out std_logic;                                        -- VRAM_ctrl_tcm_data_out_outen
			VRAM_ctrl_tcm_chipselect_n_out : out std_logic_vector(0 downto 0);                     -- VRAM_ctrl_tcm_chipselect_n_out_out
			ROM_ctrl_tcm_chipselect_n_out  : out std_logic_vector(0 downto 0);                     -- ROM_ctrl_tcm_chipselect_n_out_out
			RAM_ctrl_tcm_chipselect_n_out  : out std_logic_vector(0 downto 0);                     -- RAM_ctrl_tcm_chipselect_n_out_out
			address                        : out std_logic_vector(15 downto 0);                    -- address_out
			r_w                            : out std_logic_vector(0 downto 0);                     -- r_w_out
			data                           : out std_logic_vector(7 downto 0);                     -- data_out
			data_in                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_in
			data_outen                     : out std_logic;                                        -- data_outen
			tcs0_request                   : in  std_logic                     := 'X';             -- request
			tcs0_grant                     : out std_logic;                                        -- grant
			tcs0_address_out               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address_out
			tcs0_write_n_out               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_data_out                  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs0_data_in                   : out std_logic_vector(7 downto 0);                     -- data_in
			tcs0_data_outen                : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcs1_request                   : in  std_logic                     := 'X';             -- request
			tcs1_grant                     : out std_logic;                                        -- grant
			tcs1_address_out               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address_out
			tcs1_write_n_out               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs1_data_out                  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs1_data_in                   : out std_logic_vector(7 downto 0);                     -- data_in
			tcs1_data_outen                : in  std_logic                     := 'X';             -- data_outen
			tcs1_chipselect_n_out          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcs2_request                   : in  std_logic                     := 'X';             -- request
			tcs2_grant                     : out std_logic;                                        -- grant
			tcs2_address_out               : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address_out
			tcs2_waitrequest_in            : out std_logic_vector(0 downto 0);                     -- waitrequest_in
			tcs2_write_n_out               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs2_data_out                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs2_data_in                   : out std_logic_vector(15 downto 0);                    -- data_in
			tcs2_data_outen                : in  std_logic                     := 'X';             -- data_outen
			tcs2_chipselect_n_out          : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component proc_PIN_share;

	component proc_BRIDGE is
		port (
			clk                                : in    std_logic                     := 'X';             -- clk
			reset                              : in    std_logic                     := 'X';             -- reset
			request                            : in    std_logic                     := 'X';             -- request
			grant                              : out   std_logic;                                        -- grant
			tcs_VRAM_ctrl_tcm_data_out         : in    std_logic_vector(15 downto 0) := (others => 'X'); -- VRAM_ctrl_tcm_data_out_out
			tcs_VRAM_ctrl_tcm_data_outen       : in    std_logic                     := 'X';             -- VRAM_ctrl_tcm_data_out_outen
			tcs_VRAM_ctrl_tcm_data_in          : out   std_logic_vector(15 downto 0);                    -- VRAM_ctrl_tcm_data_out_in
			tcs_VRAM_ctrl_tcm_chipselect_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- VRAM_ctrl_tcm_chipselect_n_out_out
			tcs_VRAM_ctrl_tcm_waitrequest_in   : out   std_logic_vector(0 downto 0);                     -- VRAM_ctrl_tcm_waitrequest_in_in
			tcs_data                           : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs_data_outen                     : in    std_logic                     := 'X';             -- data_outen
			tcs_data_in                        : out   std_logic_vector(7 downto 0);                     -- data_in
			tcs_VRAM_ctrl_tcm_address_out      : in    std_logic_vector(18 downto 0) := (others => 'X'); -- VRAM_ctrl_tcm_address_out_out
			tcs_r_w                            : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- r_w_out
			tcs_RAM_ctrl_tcm_chipselect_n_out  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- RAM_ctrl_tcm_chipselect_n_out_out
			tcs_VRAM_ctrl_tcm_write_n_out      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- VRAM_ctrl_tcm_write_n_out_out
			tcs_ROM_ctrl_tcm_chipselect_n_out  : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- ROM_ctrl_tcm_chipselect_n_out_out
			tcs_address                        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- address_out
			VRAM_ctrl_tcm_data_out             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- VRAM_ctrl_tcm_data_out
			VRAM_ctrl_tcm_chipselect_n_out     : out   std_logic_vector(0 downto 0);                     -- VRAM_ctrl_tcm_chipselect_n_out
			VRAM_ctrl_tcm_waitrequest_in       : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- VRAM_ctrl_tcm_waitrequest_in
			data                               : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			VRAM_ctrl_tcm_address_out          : out   std_logic_vector(18 downto 0);                    -- VRAM_ctrl_tcm_address_out
			r_w                                : out   std_logic_vector(0 downto 0);                     -- r_w
			RAM_ctrl_tcm_chipselect_n_out      : out   std_logic_vector(0 downto 0);                     -- RAM_ctrl_tcm_chipselect_n_out
			VRAM_ctrl_tcm_write_n_out          : out   std_logic_vector(0 downto 0);                     -- VRAM_ctrl_tcm_write_n_out
			ROM_ctrl_tcm_chipselect_n_out      : out   std_logic_vector(0 downto 0);                     -- ROM_ctrl_tcm_chipselect_n_out
			address                            : out   std_logic_vector(15 downto 0)                     -- address
		);
	end component proc_BRIDGE;

	component proc_ONCHIP_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component proc_ONCHIP_mem;

	component proc_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component proc_sysid_qsys_0;

	component proc_key_input is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(19 downto 0) := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component proc_key_input;

	component proc_VRAM_ctrl is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_waitrequest_in   : in  std_logic                     := 'X';             -- waitrequest_in
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(18 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component proc_VRAM_ctrl;

	component proc_ADC_raw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(23 downto 0) := (others => 'X')  -- export
		);
	end component proc_ADC_raw;

	component proc_TRIG_int is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component proc_TRIG_int;

	component proc_ADC_ctrl is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component proc_ADC_ctrl;

	component proc_ADC_rate is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component proc_ADC_rate;

	component proc_TRIG_delay is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component proc_TRIG_delay;

	component proc_TRIG_error is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component proc_TRIG_error;

	component proc_test_input is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component proc_test_input;

	component proc_mm_interconnect_0 is
		port (
			SYSCLK_clk_clk                           : in  std_logic                     := 'X';             -- clk
			PROC_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			PROC_data_master_address                 : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			PROC_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			PROC_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			PROC_data_master_read                    : in  std_logic                     := 'X';             -- read
			PROC_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			PROC_data_master_write                   : in  std_logic                     := 'X';             -- write
			PROC_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			PROC_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			PROC_instruction_master_address          : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			PROC_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			PROC_instruction_master_read             : in  std_logic                     := 'X';             -- read
			PROC_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			PROC_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			ADC_ctrl_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			ADC_ctrl_s1_write                        : out std_logic;                                        -- write
			ADC_ctrl_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ADC_ctrl_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			ADC_ctrl_s1_chipselect                   : out std_logic;                                        -- chipselect
			ADC_rate_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			ADC_rate_s1_write                        : out std_logic;                                        -- write
			ADC_rate_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ADC_rate_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			ADC_rate_s1_chipselect                   : out std_logic;                                        -- chipselect
			ADC_raw_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			ADC_raw_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_input_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			key_input_s1_write                       : out std_logic;                                        -- write
			key_input_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_input_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			key_input_s1_chipselect                  : out std_logic;                                        -- chipselect
			ONCHIP_mem_s1_address                    : out std_logic_vector(14 downto 0);                    -- address
			ONCHIP_mem_s1_write                      : out std_logic;                                        -- write
			ONCHIP_mem_s1_readdata                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			ONCHIP_mem_s1_writedata                  : out std_logic_vector(7 downto 0);                     -- writedata
			ONCHIP_mem_s1_chipselect                 : out std_logic;                                        -- chipselect
			ONCHIP_mem_s1_clken                      : out std_logic;                                        -- clken
			PROC_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			PROC_jtag_debug_module_write             : out std_logic;                                        -- write
			PROC_jtag_debug_module_read              : out std_logic;                                        -- read
			PROC_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PROC_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			PROC_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			PROC_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			PROC_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			RAM_ctrl_uas_address                     : out std_logic_vector(15 downto 0);                    -- address
			RAM_ctrl_uas_write                       : out std_logic;                                        -- write
			RAM_ctrl_uas_read                        : out std_logic;                                        -- read
			RAM_ctrl_uas_readdata                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			RAM_ctrl_uas_writedata                   : out std_logic_vector(7 downto 0);                     -- writedata
			RAM_ctrl_uas_burstcount                  : out std_logic_vector(0 downto 0);                     -- burstcount
			RAM_ctrl_uas_byteenable                  : out std_logic_vector(0 downto 0);                     -- byteenable
			RAM_ctrl_uas_readdatavalid               : in  std_logic                     := 'X';             -- readdatavalid
			RAM_ctrl_uas_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			RAM_ctrl_uas_lock                        : out std_logic;                                        -- lock
			RAM_ctrl_uas_debugaccess                 : out std_logic;                                        -- debugaccess
			ROM_ctrl_uas_address                     : out std_logic_vector(15 downto 0);                    -- address
			ROM_ctrl_uas_write                       : out std_logic;                                        -- write
			ROM_ctrl_uas_read                        : out std_logic;                                        -- read
			ROM_ctrl_uas_readdata                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			ROM_ctrl_uas_writedata                   : out std_logic_vector(7 downto 0);                     -- writedata
			ROM_ctrl_uas_burstcount                  : out std_logic_vector(0 downto 0);                     -- burstcount
			ROM_ctrl_uas_byteenable                  : out std_logic_vector(0 downto 0);                     -- byteenable
			ROM_ctrl_uas_readdatavalid               : in  std_logic                     := 'X';             -- readdatavalid
			ROM_ctrl_uas_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			ROM_ctrl_uas_lock                        : out std_logic;                                        -- lock
			ROM_ctrl_uas_debugaccess                 : out std_logic;                                        -- debugaccess
			sysid_qsys_0_control_slave_address       : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			test_input_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			test_input_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_ctrl_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			TRIG_ctrl_s1_write                       : out std_logic;                                        -- write
			TRIG_ctrl_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_ctrl_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			TRIG_ctrl_s1_chipselect                  : out std_logic;                                        -- chipselect
			TRIG_delay_s1_address                    : out std_logic_vector(2 downto 0);                     -- address
			TRIG_delay_s1_write                      : out std_logic;                                        -- write
			TRIG_delay_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_delay_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			TRIG_delay_s1_chipselect                 : out std_logic;                                        -- chipselect
			TRIG_error_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			TRIG_error_s1_write                      : out std_logic;                                        -- write
			TRIG_error_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_error_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			TRIG_error_s1_chipselect                 : out std_logic;                                        -- chipselect
			TRIG_int_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			TRIG_int_s1_write                        : out std_logic;                                        -- write
			TRIG_int_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_int_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			TRIG_int_s1_chipselect                   : out std_logic;                                        -- chipselect
			TRIG_level_s1_address                    : out std_logic_vector(2 downto 0);                     -- address
			TRIG_level_s1_write                      : out std_logic;                                        -- write
			TRIG_level_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TRIG_level_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			TRIG_level_s1_chipselect                 : out std_logic;                                        -- chipselect
			VRAM_ctrl_uas_address                    : out std_logic_vector(18 downto 0);                    -- address
			VRAM_ctrl_uas_write                      : out std_logic;                                        -- write
			VRAM_ctrl_uas_read                       : out std_logic;                                        -- read
			VRAM_ctrl_uas_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			VRAM_ctrl_uas_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			VRAM_ctrl_uas_burstcount                 : out std_logic_vector(1 downto 0);                     -- burstcount
			VRAM_ctrl_uas_byteenable                 : out std_logic_vector(1 downto 0);                     -- byteenable
			VRAM_ctrl_uas_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			VRAM_ctrl_uas_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			VRAM_ctrl_uas_lock                       : out std_logic;                                        -- lock
			VRAM_ctrl_uas_debugaccess                : out std_logic                                         -- debugaccess
		);
	end component proc_mm_interconnect_0;

	component proc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component proc_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal proc_jtag_debug_module_reset_reset                    : std_logic;                     -- PROC:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	signal ram_ctrl_tcm_chipselect_n_out                         : std_logic;                     -- RAM_ctrl:tcm_chipselect_n_out -> PIN_share:tcs0_chipselect_n_out
	signal ram_ctrl_tcm_grant                                    : std_logic;                     -- PIN_share:tcs0_grant -> RAM_ctrl:tcm_grant
	signal ram_ctrl_tcm_data_outen                               : std_logic;                     -- RAM_ctrl:tcm_data_outen -> PIN_share:tcs0_data_outen
	signal ram_ctrl_tcm_request                                  : std_logic;                     -- RAM_ctrl:tcm_request -> PIN_share:tcs0_request
	signal ram_ctrl_tcm_data_out                                 : std_logic_vector(7 downto 0);  -- RAM_ctrl:tcm_data_out -> PIN_share:tcs0_data_out
	signal ram_ctrl_tcm_write_n_out                              : std_logic;                     -- RAM_ctrl:tcm_write_n_out -> PIN_share:tcs0_write_n_out
	signal ram_ctrl_tcm_address_out                              : std_logic_vector(15 downto 0); -- RAM_ctrl:tcm_address_out -> PIN_share:tcs0_address_out
	signal ram_ctrl_tcm_data_in                                  : std_logic_vector(7 downto 0);  -- PIN_share:tcs0_data_in -> RAM_ctrl:tcm_data_in
	signal rom_ctrl_tcm_chipselect_n_out                         : std_logic;                     -- ROM_ctrl:tcm_chipselect_n_out -> PIN_share:tcs1_chipselect_n_out
	signal rom_ctrl_tcm_grant                                    : std_logic;                     -- PIN_share:tcs1_grant -> ROM_ctrl:tcm_grant
	signal rom_ctrl_tcm_data_outen                               : std_logic;                     -- ROM_ctrl:tcm_data_outen -> PIN_share:tcs1_data_outen
	signal rom_ctrl_tcm_request                                  : std_logic;                     -- ROM_ctrl:tcm_request -> PIN_share:tcs1_request
	signal rom_ctrl_tcm_data_out                                 : std_logic_vector(7 downto 0);  -- ROM_ctrl:tcm_data_out -> PIN_share:tcs1_data_out
	signal rom_ctrl_tcm_write_n_out                              : std_logic;                     -- ROM_ctrl:tcm_write_n_out -> PIN_share:tcs1_write_n_out
	signal rom_ctrl_tcm_address_out                              : std_logic_vector(15 downto 0); -- ROM_ctrl:tcm_address_out -> PIN_share:tcs1_address_out
	signal rom_ctrl_tcm_data_in                                  : std_logic_vector(7 downto 0);  -- PIN_share:tcs1_data_in -> ROM_ctrl:tcm_data_in
	signal pin_share_tcm_vram_ctrl_tcm_data_out_outen            : std_logic;                     -- PIN_share:VRAM_ctrl_tcm_data_outen -> BRIDGE:tcs_VRAM_ctrl_tcm_data_outen
	signal pin_share_tcm_vram_ctrl_tcm_data_out_in               : std_logic_vector(15 downto 0); -- BRIDGE:tcs_VRAM_ctrl_tcm_data_in -> PIN_share:VRAM_ctrl_tcm_data_in
	signal pin_share_tcm_grant                                   : std_logic;                     -- BRIDGE:grant -> PIN_share:grant
	signal pin_share_tcm_rom_ctrl_tcm_chipselect_n_out_out       : std_logic_vector(0 downto 0);  -- PIN_share:ROM_ctrl_tcm_chipselect_n_out -> BRIDGE:tcs_ROM_ctrl_tcm_chipselect_n_out
	signal pin_share_tcm_vram_ctrl_tcm_write_n_out_out           : std_logic_vector(0 downto 0);  -- PIN_share:VRAM_ctrl_tcm_write_n_out -> BRIDGE:tcs_VRAM_ctrl_tcm_write_n_out
	signal pin_share_tcm_ram_ctrl_tcm_chipselect_n_out_out       : std_logic_vector(0 downto 0);  -- PIN_share:RAM_ctrl_tcm_chipselect_n_out -> BRIDGE:tcs_RAM_ctrl_tcm_chipselect_n_out
	signal pin_share_tcm_vram_ctrl_tcm_chipselect_n_out_out      : std_logic_vector(0 downto 0);  -- PIN_share:VRAM_ctrl_tcm_chipselect_n_out -> BRIDGE:tcs_VRAM_ctrl_tcm_chipselect_n_out
	signal pin_share_tcm_address_out                             : std_logic_vector(15 downto 0); -- PIN_share:address -> BRIDGE:tcs_address
	signal pin_share_tcm_vram_ctrl_tcm_address_out_out           : std_logic_vector(18 downto 0); -- PIN_share:VRAM_ctrl_tcm_address_out -> BRIDGE:tcs_VRAM_ctrl_tcm_address_out
	signal pin_share_tcm_data_outen                              : std_logic;                     -- PIN_share:data_outen -> BRIDGE:tcs_data_outen
	signal pin_share_tcm_r_w_out                                 : std_logic_vector(0 downto 0);  -- PIN_share:r_w -> BRIDGE:tcs_r_w
	signal pin_share_tcm_request                                 : std_logic;                     -- PIN_share:request -> BRIDGE:request
	signal pin_share_tcm_data_out                                : std_logic_vector(7 downto 0);  -- PIN_share:data -> BRIDGE:tcs_data
	signal pin_share_tcm_vram_ctrl_tcm_data_out_out              : std_logic_vector(15 downto 0); -- PIN_share:VRAM_ctrl_tcm_data_out -> BRIDGE:tcs_VRAM_ctrl_tcm_data_out
	signal pin_share_tcm_vram_ctrl_tcm_waitrequest_in_in         : std_logic_vector(0 downto 0);  -- BRIDGE:tcs_VRAM_ctrl_tcm_waitrequest_in -> PIN_share:VRAM_ctrl_tcm_waitrequest_in
	signal pin_share_tcm_data_in                                 : std_logic_vector(7 downto 0);  -- BRIDGE:tcs_data_in -> PIN_share:data_in
	signal vram_ctrl_tcm_chipselect_n_out                        : std_logic;                     -- VRAM_ctrl:tcm_chipselect_n_out -> PIN_share:tcs2_chipselect_n_out
	signal vram_ctrl_tcm_grant                                   : std_logic;                     -- PIN_share:tcs2_grant -> VRAM_ctrl:tcm_grant
	signal vram_ctrl_tcm_data_outen                              : std_logic;                     -- VRAM_ctrl:tcm_data_outen -> PIN_share:tcs2_data_outen
	signal vram_ctrl_tcm_request                                 : std_logic;                     -- VRAM_ctrl:tcm_request -> PIN_share:tcs2_request
	signal vram_ctrl_tcm_data_out                                : std_logic_vector(15 downto 0); -- VRAM_ctrl:tcm_data_out -> PIN_share:tcs2_data_out
	signal vram_ctrl_tcm_write_n_out                             : std_logic;                     -- VRAM_ctrl:tcm_write_n_out -> PIN_share:tcs2_write_n_out
	signal vram_ctrl_tcm_address_out                             : std_logic_vector(18 downto 0); -- VRAM_ctrl:tcm_address_out -> PIN_share:tcs2_address_out
	signal vram_ctrl_tcm_data_in                                 : std_logic_vector(15 downto 0); -- PIN_share:tcs2_data_in -> VRAM_ctrl:tcm_data_in
	signal vram_ctrl_tcm_waitrequest_in                          : std_logic;                     -- PIN_share:tcs2_waitrequest_in -> VRAM_ctrl:tcm_waitrequest_in
	signal mm_interconnect_0_vram_ctrl_uas_waitrequest           : std_logic;                     -- VRAM_ctrl:uas_waitrequest -> mm_interconnect_0:VRAM_ctrl_uas_waitrequest
	signal mm_interconnect_0_vram_ctrl_uas_burstcount            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VRAM_ctrl_uas_burstcount -> VRAM_ctrl:uas_burstcount
	signal mm_interconnect_0_vram_ctrl_uas_writedata             : std_logic_vector(15 downto 0); -- mm_interconnect_0:VRAM_ctrl_uas_writedata -> VRAM_ctrl:uas_writedata
	signal mm_interconnect_0_vram_ctrl_uas_address               : std_logic_vector(18 downto 0); -- mm_interconnect_0:VRAM_ctrl_uas_address -> VRAM_ctrl:uas_address
	signal mm_interconnect_0_vram_ctrl_uas_lock                  : std_logic;                     -- mm_interconnect_0:VRAM_ctrl_uas_lock -> VRAM_ctrl:uas_lock
	signal mm_interconnect_0_vram_ctrl_uas_write                 : std_logic;                     -- mm_interconnect_0:VRAM_ctrl_uas_write -> VRAM_ctrl:uas_write
	signal mm_interconnect_0_vram_ctrl_uas_read                  : std_logic;                     -- mm_interconnect_0:VRAM_ctrl_uas_read -> VRAM_ctrl:uas_read
	signal mm_interconnect_0_vram_ctrl_uas_readdata              : std_logic_vector(15 downto 0); -- VRAM_ctrl:uas_readdata -> mm_interconnect_0:VRAM_ctrl_uas_readdata
	signal mm_interconnect_0_vram_ctrl_uas_debugaccess           : std_logic;                     -- mm_interconnect_0:VRAM_ctrl_uas_debugaccess -> VRAM_ctrl:uas_debugaccess
	signal mm_interconnect_0_vram_ctrl_uas_readdatavalid         : std_logic;                     -- VRAM_ctrl:uas_readdatavalid -> mm_interconnect_0:VRAM_ctrl_uas_readdatavalid
	signal mm_interconnect_0_vram_ctrl_uas_byteenable            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VRAM_ctrl_uas_byteenable -> VRAM_ctrl:uas_byteenable
	signal mm_interconnect_0_trig_int_s1_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:TRIG_int_s1_writedata -> TRIG_int:writedata
	signal mm_interconnect_0_trig_int_s1_address                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TRIG_int_s1_address -> TRIG_int:address
	signal mm_interconnect_0_trig_int_s1_chipselect              : std_logic;                     -- mm_interconnect_0:TRIG_int_s1_chipselect -> TRIG_int:chipselect
	signal mm_interconnect_0_trig_int_s1_write                   : std_logic;                     -- mm_interconnect_0:TRIG_int_s1_write -> mm_interconnect_0_trig_int_s1_write:in
	signal mm_interconnect_0_trig_int_s1_readdata                : std_logic_vector(31 downto 0); -- TRIG_int:readdata -> mm_interconnect_0:TRIG_int_s1_readdata
	signal mm_interconnect_0_key_input_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_input_s1_writedata -> key_input:writedata
	signal mm_interconnect_0_key_input_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_input_s1_address -> key_input:address
	signal mm_interconnect_0_key_input_s1_chipselect             : std_logic;                     -- mm_interconnect_0:key_input_s1_chipselect -> key_input:chipselect
	signal mm_interconnect_0_key_input_s1_write                  : std_logic;                     -- mm_interconnect_0:key_input_s1_write -> mm_interconnect_0_key_input_s1_write:in
	signal mm_interconnect_0_key_input_s1_readdata               : std_logic_vector(31 downto 0); -- key_input:readdata -> mm_interconnect_0:key_input_s1_readdata
	signal mm_interconnect_0_ram_ctrl_uas_waitrequest            : std_logic;                     -- RAM_ctrl:uas_waitrequest -> mm_interconnect_0:RAM_ctrl_uas_waitrequest
	signal mm_interconnect_0_ram_ctrl_uas_burstcount             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:RAM_ctrl_uas_burstcount -> RAM_ctrl:uas_burstcount
	signal mm_interconnect_0_ram_ctrl_uas_writedata              : std_logic_vector(7 downto 0);  -- mm_interconnect_0:RAM_ctrl_uas_writedata -> RAM_ctrl:uas_writedata
	signal mm_interconnect_0_ram_ctrl_uas_address                : std_logic_vector(15 downto 0); -- mm_interconnect_0:RAM_ctrl_uas_address -> RAM_ctrl:uas_address
	signal mm_interconnect_0_ram_ctrl_uas_lock                   : std_logic;                     -- mm_interconnect_0:RAM_ctrl_uas_lock -> RAM_ctrl:uas_lock
	signal mm_interconnect_0_ram_ctrl_uas_write                  : std_logic;                     -- mm_interconnect_0:RAM_ctrl_uas_write -> RAM_ctrl:uas_write
	signal mm_interconnect_0_ram_ctrl_uas_read                   : std_logic;                     -- mm_interconnect_0:RAM_ctrl_uas_read -> RAM_ctrl:uas_read
	signal mm_interconnect_0_ram_ctrl_uas_readdata               : std_logic_vector(7 downto 0);  -- RAM_ctrl:uas_readdata -> mm_interconnect_0:RAM_ctrl_uas_readdata
	signal mm_interconnect_0_ram_ctrl_uas_debugaccess            : std_logic;                     -- mm_interconnect_0:RAM_ctrl_uas_debugaccess -> RAM_ctrl:uas_debugaccess
	signal mm_interconnect_0_ram_ctrl_uas_readdatavalid          : std_logic;                     -- RAM_ctrl:uas_readdatavalid -> mm_interconnect_0:RAM_ctrl_uas_readdatavalid
	signal mm_interconnect_0_ram_ctrl_uas_byteenable             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:RAM_ctrl_uas_byteenable -> RAM_ctrl:uas_byteenable
	signal mm_interconnect_0_trig_delay_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:TRIG_delay_s1_writedata -> TRIG_delay:writedata
	signal mm_interconnect_0_trig_delay_s1_address               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TRIG_delay_s1_address -> TRIG_delay:address
	signal mm_interconnect_0_trig_delay_s1_chipselect            : std_logic;                     -- mm_interconnect_0:TRIG_delay_s1_chipselect -> TRIG_delay:chipselect
	signal mm_interconnect_0_trig_delay_s1_write                 : std_logic;                     -- mm_interconnect_0:TRIG_delay_s1_write -> mm_interconnect_0_trig_delay_s1_write:in
	signal mm_interconnect_0_trig_delay_s1_readdata              : std_logic_vector(31 downto 0); -- TRIG_delay:readdata -> mm_interconnect_0:TRIG_delay_s1_readdata
	signal mm_interconnect_0_test_input_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:test_input_s1_address -> test_input:address
	signal mm_interconnect_0_test_input_s1_readdata              : std_logic_vector(31 downto 0); -- test_input:readdata -> mm_interconnect_0:test_input_s1_readdata
	signal mm_interconnect_0_rom_ctrl_uas_waitrequest            : std_logic;                     -- ROM_ctrl:uas_waitrequest -> mm_interconnect_0:ROM_ctrl_uas_waitrequest
	signal mm_interconnect_0_rom_ctrl_uas_burstcount             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ROM_ctrl_uas_burstcount -> ROM_ctrl:uas_burstcount
	signal mm_interconnect_0_rom_ctrl_uas_writedata              : std_logic_vector(7 downto 0);  -- mm_interconnect_0:ROM_ctrl_uas_writedata -> ROM_ctrl:uas_writedata
	signal mm_interconnect_0_rom_ctrl_uas_address                : std_logic_vector(15 downto 0); -- mm_interconnect_0:ROM_ctrl_uas_address -> ROM_ctrl:uas_address
	signal mm_interconnect_0_rom_ctrl_uas_lock                   : std_logic;                     -- mm_interconnect_0:ROM_ctrl_uas_lock -> ROM_ctrl:uas_lock
	signal mm_interconnect_0_rom_ctrl_uas_write                  : std_logic;                     -- mm_interconnect_0:ROM_ctrl_uas_write -> ROM_ctrl:uas_write
	signal mm_interconnect_0_rom_ctrl_uas_read                   : std_logic;                     -- mm_interconnect_0:ROM_ctrl_uas_read -> ROM_ctrl:uas_read
	signal mm_interconnect_0_rom_ctrl_uas_readdata               : std_logic_vector(7 downto 0);  -- ROM_ctrl:uas_readdata -> mm_interconnect_0:ROM_ctrl_uas_readdata
	signal mm_interconnect_0_rom_ctrl_uas_debugaccess            : std_logic;                     -- mm_interconnect_0:ROM_ctrl_uas_debugaccess -> ROM_ctrl:uas_debugaccess
	signal mm_interconnect_0_rom_ctrl_uas_readdatavalid          : std_logic;                     -- ROM_ctrl:uas_readdatavalid -> mm_interconnect_0:ROM_ctrl_uas_readdatavalid
	signal mm_interconnect_0_rom_ctrl_uas_byteenable             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ROM_ctrl_uas_byteenable -> ROM_ctrl:uas_byteenable
	signal mm_interconnect_0_proc_jtag_debug_module_waitrequest  : std_logic;                     -- PROC:jtag_debug_module_waitrequest -> mm_interconnect_0:PROC_jtag_debug_module_waitrequest
	signal mm_interconnect_0_proc_jtag_debug_module_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_0:PROC_jtag_debug_module_writedata -> PROC:jtag_debug_module_writedata
	signal mm_interconnect_0_proc_jtag_debug_module_address      : std_logic_vector(8 downto 0);  -- mm_interconnect_0:PROC_jtag_debug_module_address -> PROC:jtag_debug_module_address
	signal mm_interconnect_0_proc_jtag_debug_module_write        : std_logic;                     -- mm_interconnect_0:PROC_jtag_debug_module_write -> PROC:jtag_debug_module_write
	signal mm_interconnect_0_proc_jtag_debug_module_read         : std_logic;                     -- mm_interconnect_0:PROC_jtag_debug_module_read -> PROC:jtag_debug_module_read
	signal mm_interconnect_0_proc_jtag_debug_module_readdata     : std_logic_vector(31 downto 0); -- PROC:jtag_debug_module_readdata -> mm_interconnect_0:PROC_jtag_debug_module_readdata
	signal mm_interconnect_0_proc_jtag_debug_module_debugaccess  : std_logic;                     -- mm_interconnect_0:PROC_jtag_debug_module_debugaccess -> PROC:jtag_debug_module_debugaccess
	signal mm_interconnect_0_proc_jtag_debug_module_byteenable   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:PROC_jtag_debug_module_byteenable -> PROC:jtag_debug_module_byteenable
	signal proc_data_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:PROC_data_master_waitrequest -> PROC:d_waitrequest
	signal proc_data_master_writedata                            : std_logic_vector(31 downto 0); -- PROC:d_writedata -> mm_interconnect_0:PROC_data_master_writedata
	signal proc_data_master_address                              : std_logic_vector(20 downto 0); -- PROC:d_address -> mm_interconnect_0:PROC_data_master_address
	signal proc_data_master_write                                : std_logic;                     -- PROC:d_write -> mm_interconnect_0:PROC_data_master_write
	signal proc_data_master_read                                 : std_logic;                     -- PROC:d_read -> mm_interconnect_0:PROC_data_master_read
	signal proc_data_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:PROC_data_master_readdata -> PROC:d_readdata
	signal proc_data_master_debugaccess                          : std_logic;                     -- PROC:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:PROC_data_master_debugaccess
	signal proc_data_master_byteenable                           : std_logic_vector(3 downto 0);  -- PROC:d_byteenable -> mm_interconnect_0:PROC_data_master_byteenable
	signal mm_interconnect_0_adc_rate_s1_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ADC_rate_s1_writedata -> ADC_rate:writedata
	signal mm_interconnect_0_adc_rate_s1_address                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ADC_rate_s1_address -> ADC_rate:address
	signal mm_interconnect_0_adc_rate_s1_chipselect              : std_logic;                     -- mm_interconnect_0:ADC_rate_s1_chipselect -> ADC_rate:chipselect
	signal mm_interconnect_0_adc_rate_s1_write                   : std_logic;                     -- mm_interconnect_0:ADC_rate_s1_write -> mm_interconnect_0_adc_rate_s1_write:in
	signal mm_interconnect_0_adc_rate_s1_readdata                : std_logic_vector(31 downto 0); -- ADC_rate:readdata -> mm_interconnect_0:ADC_rate_s1_readdata
	signal mm_interconnect_0_adc_raw_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ADC_raw_s1_address -> ADC_raw:address
	signal mm_interconnect_0_adc_raw_s1_readdata                 : std_logic_vector(31 downto 0); -- ADC_raw:readdata -> mm_interconnect_0:ADC_raw_s1_readdata
	signal mm_interconnect_0_adc_ctrl_s1_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ADC_ctrl_s1_writedata -> ADC_ctrl:writedata
	signal mm_interconnect_0_adc_ctrl_s1_address                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ADC_ctrl_s1_address -> ADC_ctrl:address
	signal mm_interconnect_0_adc_ctrl_s1_chipselect              : std_logic;                     -- mm_interconnect_0:ADC_ctrl_s1_chipselect -> ADC_ctrl:chipselect
	signal mm_interconnect_0_adc_ctrl_s1_write                   : std_logic;                     -- mm_interconnect_0:ADC_ctrl_s1_write -> mm_interconnect_0_adc_ctrl_s1_write:in
	signal mm_interconnect_0_adc_ctrl_s1_readdata                : std_logic_vector(31 downto 0); -- ADC_ctrl:readdata -> mm_interconnect_0:ADC_ctrl_s1_readdata
	signal mm_interconnect_0_trig_ctrl_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:TRIG_ctrl_s1_writedata -> TRIG_ctrl:writedata
	signal mm_interconnect_0_trig_ctrl_s1_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TRIG_ctrl_s1_address -> TRIG_ctrl:address
	signal mm_interconnect_0_trig_ctrl_s1_chipselect             : std_logic;                     -- mm_interconnect_0:TRIG_ctrl_s1_chipselect -> TRIG_ctrl:chipselect
	signal mm_interconnect_0_trig_ctrl_s1_write                  : std_logic;                     -- mm_interconnect_0:TRIG_ctrl_s1_write -> mm_interconnect_0_trig_ctrl_s1_write:in
	signal mm_interconnect_0_trig_ctrl_s1_readdata               : std_logic_vector(31 downto 0); -- TRIG_ctrl:readdata -> mm_interconnect_0:TRIG_ctrl_s1_readdata
	signal mm_interconnect_0_trig_level_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:TRIG_level_s1_writedata -> TRIG_level:writedata
	signal mm_interconnect_0_trig_level_s1_address               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TRIG_level_s1_address -> TRIG_level:address
	signal mm_interconnect_0_trig_level_s1_chipselect            : std_logic;                     -- mm_interconnect_0:TRIG_level_s1_chipselect -> TRIG_level:chipselect
	signal mm_interconnect_0_trig_level_s1_write                 : std_logic;                     -- mm_interconnect_0:TRIG_level_s1_write -> mm_interconnect_0_trig_level_s1_write:in
	signal mm_interconnect_0_trig_level_s1_readdata              : std_logic_vector(31 downto 0); -- TRIG_level:readdata -> mm_interconnect_0:TRIG_level_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_writedata             : std_logic_vector(7 downto 0);  -- mm_interconnect_0:ONCHIP_mem_s1_writedata -> ONCHIP_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_address               : std_logic_vector(14 downto 0); -- mm_interconnect_0:ONCHIP_mem_s1_address -> ONCHIP_mem:address
	signal mm_interconnect_0_onchip_mem_s1_chipselect            : std_logic;                     -- mm_interconnect_0:ONCHIP_mem_s1_chipselect -> ONCHIP_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_clken                 : std_logic;                     -- mm_interconnect_0:ONCHIP_mem_s1_clken -> ONCHIP_mem:clken
	signal mm_interconnect_0_onchip_mem_s1_write                 : std_logic;                     -- mm_interconnect_0:ONCHIP_mem_s1_write -> ONCHIP_mem:write
	signal mm_interconnect_0_onchip_mem_s1_readdata              : std_logic_vector(7 downto 0);  -- ONCHIP_mem:readdata -> mm_interconnect_0:ONCHIP_mem_s1_readdata
	signal mm_interconnect_0_trig_error_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:TRIG_error_s1_writedata -> TRIG_error:writedata
	signal mm_interconnect_0_trig_error_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TRIG_error_s1_address -> TRIG_error:address
	signal mm_interconnect_0_trig_error_s1_chipselect            : std_logic;                     -- mm_interconnect_0:TRIG_error_s1_chipselect -> TRIG_error:chipselect
	signal mm_interconnect_0_trig_error_s1_write                 : std_logic;                     -- mm_interconnect_0:TRIG_error_s1_write -> mm_interconnect_0_trig_error_s1_write:in
	signal mm_interconnect_0_trig_error_s1_readdata              : std_logic_vector(31 downto 0); -- TRIG_error:readdata -> mm_interconnect_0:TRIG_error_s1_readdata
	signal proc_instruction_master_waitrequest                   : std_logic;                     -- mm_interconnect_0:PROC_instruction_master_waitrequest -> PROC:i_waitrequest
	signal proc_instruction_master_address                       : std_logic_vector(20 downto 0); -- PROC:i_address -> mm_interconnect_0:PROC_instruction_master_address
	signal proc_instruction_master_read                          : std_logic;                     -- PROC:i_read -> mm_interconnect_0:PROC_instruction_master_read
	signal proc_instruction_master_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:PROC_instruction_master_readdata -> PROC:i_readdata
	signal proc_instruction_master_readdatavalid                 : std_logic;                     -- mm_interconnect_0:PROC_instruction_master_readdatavalid -> PROC:i_readdatavalid
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal irq_mapper_receiver0_irq                              : std_logic;                     -- key_input:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                              : std_logic;                     -- TRIG_int:irq -> irq_mapper:receiver1_irq
	signal proc_d_irq_irq                                        : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> PROC:d_irq
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [BRIDGE:reset, ONCHIP_mem:reset, PIN_share:reset_reset, RAM_ctrl:reset_reset, ROM_ctrl:reset_reset, VRAM_ctrl:reset_reset, irq_mapper:reset, mm_interconnect_0:PROC_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                    : std_logic;                     -- rst_controller:reset_req -> [ONCHIP_mem:reset_req, PROC:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_trig_int_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_trig_int_s1_write:inv -> TRIG_int:write_n
	signal mm_interconnect_0_key_input_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_key_input_s1_write:inv -> key_input:write_n
	signal mm_interconnect_0_trig_delay_s1_write_ports_inv       : std_logic;                     -- mm_interconnect_0_trig_delay_s1_write:inv -> TRIG_delay:write_n
	signal mm_interconnect_0_adc_rate_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_adc_rate_s1_write:inv -> ADC_rate:write_n
	signal mm_interconnect_0_adc_ctrl_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_adc_ctrl_s1_write:inv -> ADC_ctrl:write_n
	signal mm_interconnect_0_trig_ctrl_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_trig_ctrl_s1_write:inv -> TRIG_ctrl:write_n
	signal mm_interconnect_0_trig_level_s1_write_ports_inv       : std_logic;                     -- mm_interconnect_0_trig_level_s1_write:inv -> TRIG_level:write_n
	signal mm_interconnect_0_trig_error_s1_write_ports_inv       : std_logic;                     -- mm_interconnect_0_trig_error_s1_write:inv -> TRIG_error:write_n
	signal rst_controller_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [ADC_ctrl:reset_n, ADC_rate:reset_n, ADC_raw:reset_n, PROC:reset_n, TRIG_ctrl:reset_n, TRIG_delay:reset_n, TRIG_error:reset_n, TRIG_int:reset_n, TRIG_level:reset_n, key_input:reset_n, sysid_qsys_0:reset_n, test_input:reset_n]

begin

	proc : component proc_PROC
		port map (
			clk                                   => clk_clk,                                              --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,             --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                             => proc_data_master_address,                             --               data_master.address
			d_byteenable                          => proc_data_master_byteenable,                          --                          .byteenable
			d_read                                => proc_data_master_read,                                --                          .read
			d_readdata                            => proc_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => proc_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => proc_data_master_write,                               --                          .write
			d_writedata                           => proc_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => proc_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => proc_instruction_master_address,                      --        instruction_master.address
			i_read                                => proc_instruction_master_read,                         --                          .read
			i_readdata                            => proc_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => proc_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => proc_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => proc_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => proc_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_proc_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_proc_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_proc_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_proc_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_proc_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_proc_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_proc_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_proc_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                  -- custom_instruction_master.readra
		);

	ram_ctrl : component proc_RAM_ctrl
		generic map (
			TCM_ADDRESS_W                  => 16,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 12,
			TCM_WRITE_WAIT                 => 8,
			TCM_SETUP_WAIT                 => 12,
			TCM_DATA_HOLD                  => 0,
			TCM_TURNAROUND_TIME            => 1,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_clk,                                      --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,               -- reset.reset
			uas_address          => mm_interconnect_0_ram_ctrl_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_ram_ctrl_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_ram_ctrl_uas_read,          --      .read
			uas_write            => mm_interconnect_0_ram_ctrl_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_ram_ctrl_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_ram_ctrl_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_ram_ctrl_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_ram_ctrl_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_ram_ctrl_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_ram_ctrl_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_ram_ctrl_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => ram_ctrl_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_chipselect_n_out => ram_ctrl_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => ram_ctrl_tcm_request,                         --      .request
			tcm_grant            => ram_ctrl_tcm_grant,                           --      .grant
			tcm_address_out      => ram_ctrl_tcm_address_out,                     --      .address_out
			tcm_data_out         => ram_ctrl_tcm_data_out,                        --      .data_out
			tcm_data_outen       => ram_ctrl_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => ram_ctrl_tcm_data_in                          --      .data_in
		);

	rom_ctrl : component proc_ROM_ctrl
		generic map (
			TCM_ADDRESS_W                  => 16,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 8,
			TCM_WRITE_WAIT                 => 8,
			TCM_SETUP_WAIT                 => 4,
			TCM_DATA_HOLD                  => 4,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 1,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_clk,                                      --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,               -- reset.reset
			uas_address          => mm_interconnect_0_rom_ctrl_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_rom_ctrl_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_rom_ctrl_uas_read,          --      .read
			uas_write            => mm_interconnect_0_rom_ctrl_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_rom_ctrl_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_rom_ctrl_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_rom_ctrl_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_rom_ctrl_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_rom_ctrl_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_rom_ctrl_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_rom_ctrl_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => rom_ctrl_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_chipselect_n_out => rom_ctrl_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_request          => rom_ctrl_tcm_request,                         --      .request
			tcm_grant            => rom_ctrl_tcm_grant,                           --      .grant
			tcm_address_out      => rom_ctrl_tcm_address_out,                     --      .address_out
			tcm_data_out         => rom_ctrl_tcm_data_out,                        --      .data_out
			tcm_data_outen       => rom_ctrl_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => rom_ctrl_tcm_data_in                          --      .data_in
		);

	pin_share : component proc_PIN_share
		port map (
			clk_clk                        => clk_clk,                                          --   clk.clk
			reset_reset                    => rst_controller_reset_out_reset,                   -- reset.reset
			request                        => pin_share_tcm_request,                            --   tcm.request
			grant                          => pin_share_tcm_grant,                              --      .grant
			VRAM_ctrl_tcm_address_out      => pin_share_tcm_vram_ctrl_tcm_address_out_out,      --      .VRAM_ctrl_tcm_address_out_out
			VRAM_ctrl_tcm_waitrequest_in   => pin_share_tcm_vram_ctrl_tcm_waitrequest_in_in,    --      .VRAM_ctrl_tcm_waitrequest_in_in
			VRAM_ctrl_tcm_write_n_out      => pin_share_tcm_vram_ctrl_tcm_write_n_out_out,      --      .VRAM_ctrl_tcm_write_n_out_out
			VRAM_ctrl_tcm_data_out         => pin_share_tcm_vram_ctrl_tcm_data_out_out,         --      .VRAM_ctrl_tcm_data_out_out
			VRAM_ctrl_tcm_data_in          => pin_share_tcm_vram_ctrl_tcm_data_out_in,          --      .VRAM_ctrl_tcm_data_out_in
			VRAM_ctrl_tcm_data_outen       => pin_share_tcm_vram_ctrl_tcm_data_out_outen,       --      .VRAM_ctrl_tcm_data_out_outen
			VRAM_ctrl_tcm_chipselect_n_out => pin_share_tcm_vram_ctrl_tcm_chipselect_n_out_out, --      .VRAM_ctrl_tcm_chipselect_n_out_out
			ROM_ctrl_tcm_chipselect_n_out  => pin_share_tcm_rom_ctrl_tcm_chipselect_n_out_out,  --      .ROM_ctrl_tcm_chipselect_n_out_out
			RAM_ctrl_tcm_chipselect_n_out  => pin_share_tcm_ram_ctrl_tcm_chipselect_n_out_out,  --      .RAM_ctrl_tcm_chipselect_n_out_out
			address                        => pin_share_tcm_address_out,                        --      .address_out
			r_w                            => pin_share_tcm_r_w_out,                            --      .r_w_out
			data                           => pin_share_tcm_data_out,                           --      .data_out
			data_in                        => pin_share_tcm_data_in,                            --      .data_in
			data_outen                     => pin_share_tcm_data_outen,                         --      .data_outen
			tcs0_request                   => ram_ctrl_tcm_request,                             --  tcs0.request
			tcs0_grant                     => ram_ctrl_tcm_grant,                               --      .grant
			tcs0_address_out               => ram_ctrl_tcm_address_out,                         --      .address_out
			tcs0_write_n_out(0)            => ram_ctrl_tcm_write_n_out,                         --      .write_n_out
			tcs0_data_out                  => ram_ctrl_tcm_data_out,                            --      .data_out
			tcs0_data_in                   => ram_ctrl_tcm_data_in,                             --      .data_in
			tcs0_data_outen                => ram_ctrl_tcm_data_outen,                          --      .data_outen
			tcs0_chipselect_n_out(0)       => ram_ctrl_tcm_chipselect_n_out,                    --      .chipselect_n_out
			tcs1_request                   => rom_ctrl_tcm_request,                             --  tcs1.request
			tcs1_grant                     => rom_ctrl_tcm_grant,                               --      .grant
			tcs1_address_out               => rom_ctrl_tcm_address_out,                         --      .address_out
			tcs1_write_n_out(0)            => rom_ctrl_tcm_write_n_out,                         --      .write_n_out
			tcs1_data_out                  => rom_ctrl_tcm_data_out,                            --      .data_out
			tcs1_data_in                   => rom_ctrl_tcm_data_in,                             --      .data_in
			tcs1_data_outen                => rom_ctrl_tcm_data_outen,                          --      .data_outen
			tcs1_chipselect_n_out(0)       => rom_ctrl_tcm_chipselect_n_out,                    --      .chipselect_n_out
			tcs2_request                   => vram_ctrl_tcm_request,                            --  tcs2.request
			tcs2_grant                     => vram_ctrl_tcm_grant,                              --      .grant
			tcs2_address_out               => vram_ctrl_tcm_address_out,                        --      .address_out
			tcs2_waitrequest_in(0)         => vram_ctrl_tcm_waitrequest_in,                     --      .waitrequest_in
			tcs2_write_n_out(0)            => vram_ctrl_tcm_write_n_out,                        --      .write_n_out
			tcs2_data_out                  => vram_ctrl_tcm_data_out,                           --      .data_out
			tcs2_data_in                   => vram_ctrl_tcm_data_in,                            --      .data_in
			tcs2_data_outen                => vram_ctrl_tcm_data_outen,                         --      .data_outen
			tcs2_chipselect_n_out(0)       => vram_ctrl_tcm_chipselect_n_out                    --      .chipselect_n_out
		);

	bridge : component proc_BRIDGE
		port map (
			clk                                => clk_clk,                                          --   clk.clk
			reset                              => rst_controller_reset_out_reset,                   -- reset.reset
			request                            => pin_share_tcm_request,                            --   tcs.request
			grant                              => pin_share_tcm_grant,                              --      .grant
			tcs_VRAM_ctrl_tcm_data_out         => pin_share_tcm_vram_ctrl_tcm_data_out_out,         --      .VRAM_ctrl_tcm_data_out_out
			tcs_VRAM_ctrl_tcm_data_outen       => pin_share_tcm_vram_ctrl_tcm_data_out_outen,       --      .VRAM_ctrl_tcm_data_out_outen
			tcs_VRAM_ctrl_tcm_data_in          => pin_share_tcm_vram_ctrl_tcm_data_out_in,          --      .VRAM_ctrl_tcm_data_out_in
			tcs_VRAM_ctrl_tcm_chipselect_n_out => pin_share_tcm_vram_ctrl_tcm_chipselect_n_out_out, --      .VRAM_ctrl_tcm_chipselect_n_out_out
			tcs_VRAM_ctrl_tcm_waitrequest_in   => pin_share_tcm_vram_ctrl_tcm_waitrequest_in_in,    --      .VRAM_ctrl_tcm_waitrequest_in_in
			tcs_data                           => pin_share_tcm_data_out,                           --      .data_out
			tcs_data_outen                     => pin_share_tcm_data_outen,                         --      .data_outen
			tcs_data_in                        => pin_share_tcm_data_in,                            --      .data_in
			tcs_VRAM_ctrl_tcm_address_out      => pin_share_tcm_vram_ctrl_tcm_address_out_out,      --      .VRAM_ctrl_tcm_address_out_out
			tcs_r_w                            => pin_share_tcm_r_w_out,                            --      .r_w_out
			tcs_RAM_ctrl_tcm_chipselect_n_out  => pin_share_tcm_ram_ctrl_tcm_chipselect_n_out_out,  --      .RAM_ctrl_tcm_chipselect_n_out_out
			tcs_VRAM_ctrl_tcm_write_n_out      => pin_share_tcm_vram_ctrl_tcm_write_n_out_out,      --      .VRAM_ctrl_tcm_write_n_out_out
			tcs_ROM_ctrl_tcm_chipselect_n_out  => pin_share_tcm_rom_ctrl_tcm_chipselect_n_out_out,  --      .ROM_ctrl_tcm_chipselect_n_out_out
			tcs_address                        => pin_share_tcm_address_out,                        --      .address_out
			VRAM_ctrl_tcm_data_out             => bridge_out_VRAM_ctrl_tcm_data_out,                --   out.VRAM_ctrl_tcm_data_out
			VRAM_ctrl_tcm_chipselect_n_out     => bridge_out_VRAM_ctrl_tcm_chipselect_n_out,        --      .VRAM_ctrl_tcm_chipselect_n_out
			VRAM_ctrl_tcm_waitrequest_in       => bridge_out_VRAM_ctrl_tcm_waitrequest_in,          --      .VRAM_ctrl_tcm_waitrequest_in
			data                               => bridge_out_data,                                  --      .data
			VRAM_ctrl_tcm_address_out          => bridge_out_VRAM_ctrl_tcm_address_out,             --      .VRAM_ctrl_tcm_address_out
			r_w                                => bridge_out_r_w,                                   --      .r_w
			RAM_ctrl_tcm_chipselect_n_out      => bridge_out_RAM_ctrl_tcm_chipselect_n_out,         --      .RAM_ctrl_tcm_chipselect_n_out
			VRAM_ctrl_tcm_write_n_out          => bridge_out_VRAM_ctrl_tcm_write_n_out,             --      .VRAM_ctrl_tcm_write_n_out
			ROM_ctrl_tcm_chipselect_n_out      => bridge_out_ROM_ctrl_tcm_chipselect_n_out,         --      .ROM_ctrl_tcm_chipselect_n_out
			address                            => bridge_out_address                                --      .address
		);

	onchip_mem : component proc_ONCHIP_mem
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	sysid_qsys_0 : component proc_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	key_input : component proc_key_input
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_key_input_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_input_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_input_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_input_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_input_s1_readdata,        --                    .readdata
			in_port    => key_input_export,                               -- external_connection.export
			irq        => irq_mapper_receiver0_irq                        --                 irq.irq
		);

	vram_ctrl : component proc_VRAM_ctrl
		generic map (
			TCM_ADDRESS_W                  => 19,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 0,
			TCM_WRITE_WAIT                 => 0,
			TCM_SETUP_WAIT                 => 0,
			TCM_DATA_HOLD                  => 0,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 1,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 1,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_clk,                                       --   clk.clk
			reset_reset          => rst_controller_reset_out_reset,                -- reset.reset
			uas_address          => mm_interconnect_0_vram_ctrl_uas_address,       --   uas.address
			uas_burstcount       => mm_interconnect_0_vram_ctrl_uas_burstcount,    --      .burstcount
			uas_read             => mm_interconnect_0_vram_ctrl_uas_read,          --      .read
			uas_write            => mm_interconnect_0_vram_ctrl_uas_write,         --      .write
			uas_waitrequest      => mm_interconnect_0_vram_ctrl_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid    => mm_interconnect_0_vram_ctrl_uas_readdatavalid, --      .readdatavalid
			uas_byteenable       => mm_interconnect_0_vram_ctrl_uas_byteenable,    --      .byteenable
			uas_readdata         => mm_interconnect_0_vram_ctrl_uas_readdata,      --      .readdata
			uas_writedata        => mm_interconnect_0_vram_ctrl_uas_writedata,     --      .writedata
			uas_lock             => mm_interconnect_0_vram_ctrl_uas_lock,          --      .lock
			uas_debugaccess      => mm_interconnect_0_vram_ctrl_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out      => vram_ctrl_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_chipselect_n_out => vram_ctrl_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_waitrequest_in   => vram_ctrl_tcm_waitrequest_in,                  --      .waitrequest_in
			tcm_request          => vram_ctrl_tcm_request,                         --      .request
			tcm_grant            => vram_ctrl_tcm_grant,                           --      .grant
			tcm_address_out      => vram_ctrl_tcm_address_out,                     --      .address_out
			tcm_data_out         => vram_ctrl_tcm_data_out,                        --      .data_out
			tcm_data_outen       => vram_ctrl_tcm_data_outen,                      --      .data_outen
			tcm_data_in          => vram_ctrl_tcm_data_in                          --      .data_in
		);

	adc_raw : component proc_ADC_raw
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_adc_raw_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_adc_raw_s1_readdata,    --                    .readdata
			in_port  => adc_raw_export                            -- external_connection.export
		);

	trig_int : component proc_TRIG_int
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_trig_int_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trig_int_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trig_int_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trig_int_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trig_int_s1_readdata,        --                    .readdata
			in_port    => trig_int_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                       --                 irq.irq
		);

	adc_ctrl : component proc_ADC_ctrl
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_adc_ctrl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_adc_ctrl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_adc_ctrl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_adc_ctrl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_adc_ctrl_s1_readdata,        --                    .readdata
			out_port   => adc_ctrl_export                                -- external_connection.export
		);

	adc_rate : component proc_ADC_rate
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_adc_rate_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_adc_rate_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_adc_rate_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_adc_rate_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_adc_rate_s1_readdata,        --                    .readdata
			out_port   => adc_rate_export                                -- external_connection.export
		);

	trig_ctrl : component proc_ADC_ctrl
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_trig_ctrl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trig_ctrl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trig_ctrl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trig_ctrl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trig_ctrl_s1_readdata,        --                    .readdata
			out_port   => trig_ctrl_export                                -- external_connection.export
		);

	trig_level : component proc_ADC_ctrl
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_trig_level_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trig_level_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trig_level_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trig_level_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trig_level_s1_readdata,        --                    .readdata
			out_port   => trig_level_export                                -- external_connection.export
		);

	trig_delay : component proc_TRIG_delay
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_trig_delay_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trig_delay_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trig_delay_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trig_delay_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trig_delay_s1_readdata,        --                    .readdata
			out_port   => trig_delay_export                                -- external_connection.export
		);

	trig_error : component proc_TRIG_error
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_trig_error_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_trig_error_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_trig_error_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_trig_error_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_trig_error_s1_readdata,        --                    .readdata
			out_port   => trig_errorr_export                               -- external_connection.export
		);

	test_input : component proc_test_input
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_test_input_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_test_input_s1_readdata, --                    .readdata
			in_port  => test_inp_export                           -- external_connection.export
		);

	mm_interconnect_0 : component proc_mm_interconnect_0
		port map (
			SYSCLK_clk_clk                           => clk_clk,                                               --                         SYSCLK_clk.clk
			PROC_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                        -- PROC_reset_n_reset_bridge_in_reset.reset
			PROC_data_master_address                 => proc_data_master_address,                              --                   PROC_data_master.address
			PROC_data_master_waitrequest             => proc_data_master_waitrequest,                          --                                   .waitrequest
			PROC_data_master_byteenable              => proc_data_master_byteenable,                           --                                   .byteenable
			PROC_data_master_read                    => proc_data_master_read,                                 --                                   .read
			PROC_data_master_readdata                => proc_data_master_readdata,                             --                                   .readdata
			PROC_data_master_write                   => proc_data_master_write,                                --                                   .write
			PROC_data_master_writedata               => proc_data_master_writedata,                            --                                   .writedata
			PROC_data_master_debugaccess             => proc_data_master_debugaccess,                          --                                   .debugaccess
			PROC_instruction_master_address          => proc_instruction_master_address,                       --            PROC_instruction_master.address
			PROC_instruction_master_waitrequest      => proc_instruction_master_waitrequest,                   --                                   .waitrequest
			PROC_instruction_master_read             => proc_instruction_master_read,                          --                                   .read
			PROC_instruction_master_readdata         => proc_instruction_master_readdata,                      --                                   .readdata
			PROC_instruction_master_readdatavalid    => proc_instruction_master_readdatavalid,                 --                                   .readdatavalid
			ADC_ctrl_s1_address                      => mm_interconnect_0_adc_ctrl_s1_address,                 --                        ADC_ctrl_s1.address
			ADC_ctrl_s1_write                        => mm_interconnect_0_adc_ctrl_s1_write,                   --                                   .write
			ADC_ctrl_s1_readdata                     => mm_interconnect_0_adc_ctrl_s1_readdata,                --                                   .readdata
			ADC_ctrl_s1_writedata                    => mm_interconnect_0_adc_ctrl_s1_writedata,               --                                   .writedata
			ADC_ctrl_s1_chipselect                   => mm_interconnect_0_adc_ctrl_s1_chipselect,              --                                   .chipselect
			ADC_rate_s1_address                      => mm_interconnect_0_adc_rate_s1_address,                 --                        ADC_rate_s1.address
			ADC_rate_s1_write                        => mm_interconnect_0_adc_rate_s1_write,                   --                                   .write
			ADC_rate_s1_readdata                     => mm_interconnect_0_adc_rate_s1_readdata,                --                                   .readdata
			ADC_rate_s1_writedata                    => mm_interconnect_0_adc_rate_s1_writedata,               --                                   .writedata
			ADC_rate_s1_chipselect                   => mm_interconnect_0_adc_rate_s1_chipselect,              --                                   .chipselect
			ADC_raw_s1_address                       => mm_interconnect_0_adc_raw_s1_address,                  --                         ADC_raw_s1.address
			ADC_raw_s1_readdata                      => mm_interconnect_0_adc_raw_s1_readdata,                 --                                   .readdata
			key_input_s1_address                     => mm_interconnect_0_key_input_s1_address,                --                       key_input_s1.address
			key_input_s1_write                       => mm_interconnect_0_key_input_s1_write,                  --                                   .write
			key_input_s1_readdata                    => mm_interconnect_0_key_input_s1_readdata,               --                                   .readdata
			key_input_s1_writedata                   => mm_interconnect_0_key_input_s1_writedata,              --                                   .writedata
			key_input_s1_chipselect                  => mm_interconnect_0_key_input_s1_chipselect,             --                                   .chipselect
			ONCHIP_mem_s1_address                    => mm_interconnect_0_onchip_mem_s1_address,               --                      ONCHIP_mem_s1.address
			ONCHIP_mem_s1_write                      => mm_interconnect_0_onchip_mem_s1_write,                 --                                   .write
			ONCHIP_mem_s1_readdata                   => mm_interconnect_0_onchip_mem_s1_readdata,              --                                   .readdata
			ONCHIP_mem_s1_writedata                  => mm_interconnect_0_onchip_mem_s1_writedata,             --                                   .writedata
			ONCHIP_mem_s1_chipselect                 => mm_interconnect_0_onchip_mem_s1_chipselect,            --                                   .chipselect
			ONCHIP_mem_s1_clken                      => mm_interconnect_0_onchip_mem_s1_clken,                 --                                   .clken
			PROC_jtag_debug_module_address           => mm_interconnect_0_proc_jtag_debug_module_address,      --             PROC_jtag_debug_module.address
			PROC_jtag_debug_module_write             => mm_interconnect_0_proc_jtag_debug_module_write,        --                                   .write
			PROC_jtag_debug_module_read              => mm_interconnect_0_proc_jtag_debug_module_read,         --                                   .read
			PROC_jtag_debug_module_readdata          => mm_interconnect_0_proc_jtag_debug_module_readdata,     --                                   .readdata
			PROC_jtag_debug_module_writedata         => mm_interconnect_0_proc_jtag_debug_module_writedata,    --                                   .writedata
			PROC_jtag_debug_module_byteenable        => mm_interconnect_0_proc_jtag_debug_module_byteenable,   --                                   .byteenable
			PROC_jtag_debug_module_waitrequest       => mm_interconnect_0_proc_jtag_debug_module_waitrequest,  --                                   .waitrequest
			PROC_jtag_debug_module_debugaccess       => mm_interconnect_0_proc_jtag_debug_module_debugaccess,  --                                   .debugaccess
			RAM_ctrl_uas_address                     => mm_interconnect_0_ram_ctrl_uas_address,                --                       RAM_ctrl_uas.address
			RAM_ctrl_uas_write                       => mm_interconnect_0_ram_ctrl_uas_write,                  --                                   .write
			RAM_ctrl_uas_read                        => mm_interconnect_0_ram_ctrl_uas_read,                   --                                   .read
			RAM_ctrl_uas_readdata                    => mm_interconnect_0_ram_ctrl_uas_readdata,               --                                   .readdata
			RAM_ctrl_uas_writedata                   => mm_interconnect_0_ram_ctrl_uas_writedata,              --                                   .writedata
			RAM_ctrl_uas_burstcount                  => mm_interconnect_0_ram_ctrl_uas_burstcount,             --                                   .burstcount
			RAM_ctrl_uas_byteenable                  => mm_interconnect_0_ram_ctrl_uas_byteenable,             --                                   .byteenable
			RAM_ctrl_uas_readdatavalid               => mm_interconnect_0_ram_ctrl_uas_readdatavalid,          --                                   .readdatavalid
			RAM_ctrl_uas_waitrequest                 => mm_interconnect_0_ram_ctrl_uas_waitrequest,            --                                   .waitrequest
			RAM_ctrl_uas_lock                        => mm_interconnect_0_ram_ctrl_uas_lock,                   --                                   .lock
			RAM_ctrl_uas_debugaccess                 => mm_interconnect_0_ram_ctrl_uas_debugaccess,            --                                   .debugaccess
			ROM_ctrl_uas_address                     => mm_interconnect_0_rom_ctrl_uas_address,                --                       ROM_ctrl_uas.address
			ROM_ctrl_uas_write                       => mm_interconnect_0_rom_ctrl_uas_write,                  --                                   .write
			ROM_ctrl_uas_read                        => mm_interconnect_0_rom_ctrl_uas_read,                   --                                   .read
			ROM_ctrl_uas_readdata                    => mm_interconnect_0_rom_ctrl_uas_readdata,               --                                   .readdata
			ROM_ctrl_uas_writedata                   => mm_interconnect_0_rom_ctrl_uas_writedata,              --                                   .writedata
			ROM_ctrl_uas_burstcount                  => mm_interconnect_0_rom_ctrl_uas_burstcount,             --                                   .burstcount
			ROM_ctrl_uas_byteenable                  => mm_interconnect_0_rom_ctrl_uas_byteenable,             --                                   .byteenable
			ROM_ctrl_uas_readdatavalid               => mm_interconnect_0_rom_ctrl_uas_readdatavalid,          --                                   .readdatavalid
			ROM_ctrl_uas_waitrequest                 => mm_interconnect_0_rom_ctrl_uas_waitrequest,            --                                   .waitrequest
			ROM_ctrl_uas_lock                        => mm_interconnect_0_rom_ctrl_uas_lock,                   --                                   .lock
			ROM_ctrl_uas_debugaccess                 => mm_interconnect_0_rom_ctrl_uas_debugaccess,            --                                   .debugaccess
			sysid_qsys_0_control_slave_address       => mm_interconnect_0_sysid_qsys_0_control_slave_address,  --         sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata      => mm_interconnect_0_sysid_qsys_0_control_slave_readdata, --                                   .readdata
			test_input_s1_address                    => mm_interconnect_0_test_input_s1_address,               --                      test_input_s1.address
			test_input_s1_readdata                   => mm_interconnect_0_test_input_s1_readdata,              --                                   .readdata
			TRIG_ctrl_s1_address                     => mm_interconnect_0_trig_ctrl_s1_address,                --                       TRIG_ctrl_s1.address
			TRIG_ctrl_s1_write                       => mm_interconnect_0_trig_ctrl_s1_write,                  --                                   .write
			TRIG_ctrl_s1_readdata                    => mm_interconnect_0_trig_ctrl_s1_readdata,               --                                   .readdata
			TRIG_ctrl_s1_writedata                   => mm_interconnect_0_trig_ctrl_s1_writedata,              --                                   .writedata
			TRIG_ctrl_s1_chipselect                  => mm_interconnect_0_trig_ctrl_s1_chipselect,             --                                   .chipselect
			TRIG_delay_s1_address                    => mm_interconnect_0_trig_delay_s1_address,               --                      TRIG_delay_s1.address
			TRIG_delay_s1_write                      => mm_interconnect_0_trig_delay_s1_write,                 --                                   .write
			TRIG_delay_s1_readdata                   => mm_interconnect_0_trig_delay_s1_readdata,              --                                   .readdata
			TRIG_delay_s1_writedata                  => mm_interconnect_0_trig_delay_s1_writedata,             --                                   .writedata
			TRIG_delay_s1_chipselect                 => mm_interconnect_0_trig_delay_s1_chipselect,            --                                   .chipselect
			TRIG_error_s1_address                    => mm_interconnect_0_trig_error_s1_address,               --                      TRIG_error_s1.address
			TRIG_error_s1_write                      => mm_interconnect_0_trig_error_s1_write,                 --                                   .write
			TRIG_error_s1_readdata                   => mm_interconnect_0_trig_error_s1_readdata,              --                                   .readdata
			TRIG_error_s1_writedata                  => mm_interconnect_0_trig_error_s1_writedata,             --                                   .writedata
			TRIG_error_s1_chipselect                 => mm_interconnect_0_trig_error_s1_chipselect,            --                                   .chipselect
			TRIG_int_s1_address                      => mm_interconnect_0_trig_int_s1_address,                 --                        TRIG_int_s1.address
			TRIG_int_s1_write                        => mm_interconnect_0_trig_int_s1_write,                   --                                   .write
			TRIG_int_s1_readdata                     => mm_interconnect_0_trig_int_s1_readdata,                --                                   .readdata
			TRIG_int_s1_writedata                    => mm_interconnect_0_trig_int_s1_writedata,               --                                   .writedata
			TRIG_int_s1_chipselect                   => mm_interconnect_0_trig_int_s1_chipselect,              --                                   .chipselect
			TRIG_level_s1_address                    => mm_interconnect_0_trig_level_s1_address,               --                      TRIG_level_s1.address
			TRIG_level_s1_write                      => mm_interconnect_0_trig_level_s1_write,                 --                                   .write
			TRIG_level_s1_readdata                   => mm_interconnect_0_trig_level_s1_readdata,              --                                   .readdata
			TRIG_level_s1_writedata                  => mm_interconnect_0_trig_level_s1_writedata,             --                                   .writedata
			TRIG_level_s1_chipselect                 => mm_interconnect_0_trig_level_s1_chipselect,            --                                   .chipselect
			VRAM_ctrl_uas_address                    => mm_interconnect_0_vram_ctrl_uas_address,               --                      VRAM_ctrl_uas.address
			VRAM_ctrl_uas_write                      => mm_interconnect_0_vram_ctrl_uas_write,                 --                                   .write
			VRAM_ctrl_uas_read                       => mm_interconnect_0_vram_ctrl_uas_read,                  --                                   .read
			VRAM_ctrl_uas_readdata                   => mm_interconnect_0_vram_ctrl_uas_readdata,              --                                   .readdata
			VRAM_ctrl_uas_writedata                  => mm_interconnect_0_vram_ctrl_uas_writedata,             --                                   .writedata
			VRAM_ctrl_uas_burstcount                 => mm_interconnect_0_vram_ctrl_uas_burstcount,            --                                   .burstcount
			VRAM_ctrl_uas_byteenable                 => mm_interconnect_0_vram_ctrl_uas_byteenable,            --                                   .byteenable
			VRAM_ctrl_uas_readdatavalid              => mm_interconnect_0_vram_ctrl_uas_readdatavalid,         --                                   .readdatavalid
			VRAM_ctrl_uas_waitrequest                => mm_interconnect_0_vram_ctrl_uas_waitrequest,           --                                   .waitrequest
			VRAM_ctrl_uas_lock                       => mm_interconnect_0_vram_ctrl_uas_lock,                  --                                   .lock
			VRAM_ctrl_uas_debugaccess                => mm_interconnect_0_vram_ctrl_uas_debugaccess            --                                   .debugaccess
		);

	irq_mapper : component proc_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => proc_d_irq_irq                  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => proc_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1      => proc_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_trig_int_s1_write_ports_inv <= not mm_interconnect_0_trig_int_s1_write;

	mm_interconnect_0_key_input_s1_write_ports_inv <= not mm_interconnect_0_key_input_s1_write;

	mm_interconnect_0_trig_delay_s1_write_ports_inv <= not mm_interconnect_0_trig_delay_s1_write;

	mm_interconnect_0_adc_rate_s1_write_ports_inv <= not mm_interconnect_0_adc_rate_s1_write;

	mm_interconnect_0_adc_ctrl_s1_write_ports_inv <= not mm_interconnect_0_adc_ctrl_s1_write;

	mm_interconnect_0_trig_ctrl_s1_write_ports_inv <= not mm_interconnect_0_trig_ctrl_s1_write;

	mm_interconnect_0_trig_level_s1_write_ports_inv <= not mm_interconnect_0_trig_level_s1_write;

	mm_interconnect_0_trig_error_s1_write_ports_inv <= not mm_interconnect_0_trig_error_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of proc
